// Code your design here
`include "light_package.sv"
`include "traffic_light_controller_part2_starter.sv"