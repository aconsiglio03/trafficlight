// Code your testbench here
// or browse Examples
`include "lab3_part2_tb_file.sv"